-------------------------------------------------------------------------------
-- Declaration
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package util_p is

  function is_metavalue (v : unsigned) return boolean;

end package util_p;

-------------------------------------------------------------------------------
-- Definition
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package body util_p is

  function is_metavalue (
    v : unsigned)
    return boolean is
  begin
    for i in v'range loop
      if v(i) /= '0' and v(i) /= '1' then
        return true;
      end if;
      return false;
    end loop;
  end function is_metavalue;

end package body util_p;
